library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

--This component receives the real value of the tip of the vector. Then, for every bit value, it checks if it should be painted or not according to the real value.

entity memory_writer is
	generic(ROWS : integer := 350; COLUMNS : integer := 350; BITS : integer := 32);
	port(
		clk : in std_logic := '0';
		enable : in std_logic := '0';
		rst : in std_logic := '0';
		pixel_x : out std_logic_vector(9 downto 0) := (others => '0');
		pixel_y : out std_logic_vector(9 downto 0) := (others => '0');
		pixel_on : out std_logic_vector(0 downto 0) := (others => '0')
	);

end entity;


architecture memory_writer_arq of memory_writer is
	constant AXIS_X_BIT : std_logic_vector(9 downto 0) := std_logic_vector(shift_right(to_unsigned(COLUMNS,10),1));
	constant AXIS_Y_BIT : std_logic_vector(9 downto 0) := std_logic_vector(shift_right(to_unsigned(ROWS,10),1));

	constant ONE : unsigned(BITS - 1 downto 0) := "00000000000000010000000000000000"; --1.0
	constant PIXEL_COEF : unsigned(BITS - 1 downto 0) := "00000000101011110000000000000000"; --350/2 to account for the displacement by 1

	constant POINTS_LENGTH : integer := 176;

	constant ROTATION_ANGLE : std_logic_vector(31 downto 0) := "00000000000000001011010000000000"; --0.703125 degrees

	signal unrotated_x : std_logic_vector(31 downto 0) := (others => '0');
	signal unrotated_y : std_logic_vector(31 downto 0) := (others => '0');
	
	signal cordic_to_writer_x : std_logic_vector(31 downto 0) := (others => '0');
	signal cordic_to_writer_y : std_logic_vector(31 downto 0) := (others => '0');

	signal rotation_angle_signal : std_logic_vector(31 downto 0) := (others => '0');

	component cordic is
    generic(TOTAL_BITS: integer := 32; STEPS: integer := 16);
    port(
      x_in: in std_logic_vector(TOTAL_BITS - 1 downto 0) := (others => '0');
      y_in: in std_logic_vector(TOTAL_BITS - 1 downto 0) := (others => '0');
      angle: in std_logic_vector(TOTAL_BITS - 1 downto 0) := (others => '0');
      x_out: out std_logic_vector(TOTAL_BITS - 1 downto 0) := (others => '0');
      y_out: out std_logic_vector(TOTAL_BITS - 1 downto 0) := (others => '0')
    );
  end component;

begin

	cordic_0 : cordic
    port map(
      x_in => unrotated_x,
      y_in => unrotated_y,
      angle => rotation_angle_signal,
      x_out => cordic_to_writer_x,
      y_out => cordic_to_writer_y
    );

  rotation_angle_signal <= ROTATION_ANGLE;

	
	process(clk, rst)

		variable real_x : std_logic_vector(BITS - 1 downto 0) := (others => '0');
		variable real_y : std_logic_vector(BITS - 1 downto 0) := (others => '0');

		variable moved_x : unsigned(BITS - 1 downto 0) := (others => '0');
		variable moved_y : unsigned(BITS - 1 downto 0) := (others => '0');

		variable extended_moved_x_bit : std_logic_vector(BITS * 2 - 1 downto 0) := (others => '0');
		
		variable extended_moved_y_bit_unsigned : unsigned(BITS * 2 - 1 downto 0) := (others => '0');
		variable truncated_extended_moved_y_bit_unsigned : unsigned(9 downto 0) := (others => '0');
		variable inverted_y_bit : unsigned(9 downto 0) := (others => '0');
		
		variable extended_moved_y_bit : std_logic_vector(BITS * 2 - 1 downto 0) := (others => '0');

		variable moved_x_bit : std_logic_vector(9 downto 0) := (others => '0');
		variable moved_y_bit : std_logic_vector(9 downto 0) := (others => '0');

		variable point_position : integer := 0;

		type real_point is record
			x : std_logic_vector(BITS - 1 downto 0);
			y : std_logic_vector(BITS - 1 downto 0);
		end record;
		--  The patterns to apply.
		type on_points_array is array (natural range <>) of real_point;

		variable points_to_draw : on_points_array(0 to 175) := (
					("00000000000000000000000000000000","00000000000000000000000000000000"),
					("00000000000000000000000101110110","00000000000000000000000000000000"),
					("00000000000000000000001011101100","00000000000000000000000000000000"),
					("00000000000000000000010001100011","00000000000000000000000000000000"),
					("00000000000000000000010111011001","00000000000000000000000000000000"),
					("00000000000000000000011101010000","00000000000000000000000000000000"),
					("00000000000000000000100011000110","00000000000000000000000000000000"),
					("00000000000000000000101000111101","00000000000000000000000000000000"),
					("00000000000000000000101110110011","00000000000000000000000000000000"),
					("00000000000000000000110100101010","00000000000000000000000000000000"),
					("00000000000000000000111010100000","00000000000000000000000000000000"),
					("00000000000000000001000000010111","00000000000000000000000000000000"),
					("00000000000000000001000110001101","00000000000000000000000000000000"),
					("00000000000000000001001100000100","00000000000000000000000000000000"),
					("00000000000000000001010001111010","00000000000000000000000000000000"),
					("00000000000000000001010111110001","00000000000000000000000000000000"),
					("00000000000000000001011101100111","00000000000000000000000000000000"),
					("00000000000000000001100011011110","00000000000000000000000000000000"),
					("00000000000000000001101001010100","00000000000000000000000000000000"),
					("00000000000000000001101111001011","00000000000000000000000000000000"),
					("00000000000000000001110101000001","00000000000000000000000000000000"),
					("00000000000000000001111010111000","00000000000000000000000000000000"),
					("00000000000000000010000000101110","00000000000000000000000000000000"),
					("00000000000000000010000110100101","00000000000000000000000000000000"),
					("00000000000000000010001100011011","00000000000000000000000000000000"),
					("00000000000000000010010010010010","00000000000000000000000000000000"),
					("00000000000000000010011000001000","00000000000000000000000000000000"),
					("00000000000000000010011101111111","00000000000000000000000000000000"),
					("00000000000000000010100011110101","00000000000000000000000000000000"),
					("00000000000000000010101001101100","00000000000000000000000000000000"),
					("00000000000000000010101111100010","00000000000000000000000000000000"),
					("00000000000000000010110101011001","00000000000000000000000000000000"),
					("00000000000000000010111011001111","00000000000000000000000000000000"),
					("00000000000000000011000001000110","00000000000000000000000000000000"),
					("00000000000000000011000110111100","00000000000000000000000000000000"),
					("00000000000000000011001100110011","00000000000000000000000000000000"),
					("00000000000000000011010010101001","00000000000000000000000000000000"),
					("00000000000000000011011000100000","00000000000000000000000000000000"),
					("00000000000000000011011110010110","00000000000000000000000000000000"),
					("00000000000000000011100100001101","00000000000000000000000000000000"),
					("00000000000000000011101010000011","00000000000000000000000000000000"),
					("00000000000000000011101111111010","00000000000000000000000000000000"),
					("00000000000000000011110101110000","00000000000000000000000000000000"),
					("00000000000000000011111011100111","00000000000000000000000000000000"),
					("00000000000000000100000001011101","00000000000000000000000000000000"),
					("00000000000000000100000111010100","00000000000000000000000000000000"),
					("00000000000000000100001101001010","00000000000000000000000000000000"),
					("00000000000000000100010011000001","00000000000000000000000000000000"),
					("00000000000000000100011000110111","00000000000000000000000000000000"),
					("00000000000000000100011110101110","00000000000000000000000000000000"),
					("00000000000000000100100100100100","00000000000000000000000000000000"),
					("00000000000000000100101010011011","00000000000000000000000000000000"),
					("00000000000000000100110000010001","00000000000000000000000000000000"),
					("00000000000000000100110110001000","00000000000000000000000000000000"),
					("00000000000000000100111011111110","00000000000000000000000000000000"),
					("00000000000000000101000001110101","00000000000000000000000000000000"),
					("00000000000000000101000111101011","00000000000000000000000000000000"),
					("00000000000000000101001101100010","00000000000000000000000000000000"),
					("00000000000000000101010011011000","00000000000000000000000000000000"),
					("00000000000000000101011001001110","00000000000000000000000000000000"),
					("00000000000000000101011111000101","00000000000000000000000000000000"),
					("00000000000000000101100100111011","00000000000000000000000000000000"),
					("00000000000000000101101010110010","00000000000000000000000000000000"),
					("00000000000000000101110000101000","00000000000000000000000000000000"),
					("00000000000000000101110110011111","00000000000000000000000000000000"),
					("00000000000000000101111100010101","00000000000000000000000000000000"),
					("00000000000000000110000010001100","00000000000000000000000000000000"),
					("00000000000000000110001000000010","00000000000000000000000000000000"),
					("00000000000000000110001101111001","00000000000000000000000000000000"),
					("00000000000000000110010011101111","00000000000000000000000000000000"),
					("00000000000000000110011001100110","00000000000000000000000000000000"),
					("00000000000000000110011111011100","00000000000000000000000000000000"),
					("00000000000000000110100101010011","00000000000000000000000000000000"),
					("00000000000000000110101011001001","00000000000000000000000000000000"),
					("00000000000000000110110001000000","00000000000000000000000000000000"),
					("00000000000000000110110110110110","00000000000000000000000000000000"),
					("00000000000000000110111100101101","00000000000000000000000000000000"),
					("00000000000000000111000010100011","00000000000000000000000000000000"),
					("00000000000000000111001000011010","00000000000000000000000000000000"),
					("00000000000000000111001110010000","00000000000000000000000000000000"),
					("00000000000000000111010100000111","00000000000000000000000000000000"),
					("00000000000000000111011001111101","00000000000000000000000000000000"),
					("00000000000000000111011111110100","00000000000000000000000000000000"),
					("00000000000000000111100101101010","00000000000000000000000000000000"),
					("00000000000000000111101011100001","00000000000000000000000000000000"),
					("00000000000000000111110001010111","00000000000000000000000000000000"),
					("00000000000000000111110111001110","00000000000000000000000000000000"),
					("00000000000000000111111101000100","00000000000000000000000000000000"),
					("00000000000000001000000010111011","00000000000000000000000000000000"),
					("00000000000000001000001000110001","00000000000000000000000000000000"),
					("00000000000000001000001110101000","00000000000000000000000000000000"),
					("00000000000000001000010100011110","00000000000000000000000000000000"),
					("00000000000000001000011010010101","00000000000000000000000000000000"),
					("00000000000000001000100000001011","00000000000000000000000000000000"),
					("00000000000000001000100110000010","00000000000000000000000000000000"),
					("00000000000000001000101011111000","00000000000000000000000000000000"),
					("00000000000000001000110001101111","00000000000000000000000000000000"),
					("00000000000000001000110111100101","00000000000000000000000000000000"),
					("00000000000000001000111101011100","00000000000000000000000000000000"),
					("00000000000000001001000011010010","00000000000000000000000000000000"),
					("00000000000000001001001001001001","00000000000000000000000000000000"),
					("00000000000000001001001110111111","00000000000000000000000000000000"),
					("00000000000000001001010100110110","00000000000000000000000000000000"),
					("00000000000000001001011010101100","00000000000000000000000000000000"),
					("00000000000000001001100000100011","00000000000000000000000000000000"),
					("00000000000000001001100110011001","00000000000000000000000000000000"),
					("00000000000000001001101100010000","00000000000000000000000000000000"),
					("00000000000000001001110010000110","00000000000000000000000000000000"),
					("00000000000000001001110111111101","00000000000000000000000000000000"),
					("00000000000000001001111101110011","00000000000000000000000000000000"),
					("00000000000000001010000011101010","00000000000000000000000000000000"),
					("00000000000000001010001001100000","00000000000000000000000000000000"),
					("00000000000000001010001111010111","00000000000000000000000000000000"),
					("00000000000000001010010101001101","00000000000000000000000000000000"),
					("00000000000000001010011011000100","00000000000000000000000000000000"),
					("00000000000000001010100000111010","00000000000000000000000000000000"),
					("00000000000000001010100110110001","00000000000000000000000000000000"),
					("00000000000000001010101100100111","00000000000000000000000000000000"),
					("00000000000000001010110010011101","00000000000000000000000000000000"),
					("00000000000000001010111000010100","00000000000000000000000000000000"),
					("00000000000000001010111110001010","00000000000000000000000000000000"),
					("00000000000000001011000100000001","00000000000000000000000000000000"),
					("00000000000000001011001001110111","00000000000000000000000000000000"),
					("00000000000000001011001111101110","00000000000000000000000000000000"),
					("00000000000000001011010101100100","00000000000000000000000000000000"),
					("00000000000000001011011011011011","00000000000000000000000000000000"),
					("00000000000000001011100001010001","00000000000000000000000000000000"),
					("00000000000000001011100111001000","00000000000000000000000000000000"),
					("00000000000000001011101100111110","00000000000000000000000000000000"),
					("00000000000000001011110010110101","00000000000000000000000000000000"),
					("00000000000000001011111000101011","00000000000000000000000000000000"),
					("00000000000000001011111110100010","00000000000000000000000000000000"),
					("00000000000000001100000100011000","00000000000000000000000000000000"),
					("00000000000000001100001010001111","00000000000000000000000000000000"),
					("00000000000000001100010000000101","00000000000000000000000000000000"),
					("00000000000000001100010101111100","00000000000000000000000000000000"),
					("00000000000000001100011011110010","00000000000000000000000000000000"),
					("00000000000000001100100001101001","00000000000000000000000000000000"),
					("00000000000000001100100111011111","00000000000000000000000000000000"),
					("00000000000000001100101101010110","00000000000000000000000000000000"),
					("00000000000000001100110011001100","00000000000000000000000000000000"),
					("00000000000000001100111001000011","00000000000000000000000000000000"),
					("00000000000000001100111110111001","00000000000000000000000000000000"),
					("00000000000000001101000100110000","00000000000000000000000000000000"),
					("00000000000000001101001010100110","00000000000000000000000000000000"),
					("00000000000000001101010000011101","00000000000000000000000000000000"),
					("00000000000000001101010110010011","00000000000000000000000000000000"),
					("00000000000000001101011100001010","00000000000000000000000000000000"),
					("00000000000000001101100010000000","00000000000000000000000000000000"),
					("00000000000000001101100111110111","00000000000000000000000000000000"),
					("00000000000000001101101101101101","00000000000000000000000000000000"),
					("00000000000000001101110011100100","00000000000000000000000000000000"),
					("00000000000000001101111001011010","00000000000000000000000000000000"),
					("00000000000000001101111111010001","00000000000000000000000000000000"),
					("00000000000000001110000101000111","00000000000000000000000000000000"),
					("00000000000000001110001010111110","00000000000000000000000000000000"),
					("00000000000000001110010000110100","00000000000000000000000000000000"),
					("00000000000000001110010110101011","00000000000000000000000000000000"),
					("00000000000000001110011100100001","00000000000000000000000000000000"),
					("00000000000000001110100010011000","00000000000000000000000000000000"),
					("00000000000000001110101000001110","00000000000000000000000000000000"),
					("00000000000000001110101110000101","00000000000000000000000000000000"),
					("00000000000000001110110011111011","00000000000000000000000000000000"),
					("00000000000000001110111001110010","00000000000000000000000000000000"),
					("00000000000000001110111111101000","00000000000000000000000000000000"),
					("00000000000000001111000101011111","00000000000000000000000000000000"),
					("00000000000000001111001011010101","00000000000000000000000000000000"),
					("00000000000000001111010001001100","00000000000000000000000000000000"),
					("00000000000000001111010111000010","00000000000000000000000000000000"),
					("00000000000000001111011100111001","00000000000000000000000000000000"),
					("00000000000000001111100010101111","00000000000000000000000000000000"),
					("00000000000000001111101000100110","00000000000000000000000000000000"),
					("00000000000000001111101110011100","00000000000000000000000000000000"),
					("00000000000000001111110100010011","00000000000000000000000000000000"),
					("00000000000000001111111010001001","00000000000000000000000000000000"),
					("00000000000000010000000000000000","00000000000000000000000000000000")
			);

			variable rotated_points : on_points_array(0 to 175);
	

	begin

		if(rising_edge(rst)) then --reset values
			point_position := 0;
			pixel_on <= (others => '0');
		end if;
		if(rising_edge(clk)) then

			if(enable = '1') then

				if(point_position < POINTS_LENGTH) then

					--To give time to the cordic to process the data, we shall draw the previous point and in the end set the next point to be processed
					moved_x := unsigned(points_to_draw(point_position).x) + ONE; --Move the x value to the right so that all it's posible locations are a positive number
					moved_y := unsigned(points_to_draw(point_position).y) + ONE; --Move the y value up so that all it's possible locations are a positive number

					extended_moved_x_bit := std_logic_vector(moved_x * PIXEL_COEF); --Compute the pixel location
					moved_x_bit := extended_moved_x_bit(32 + 9 downto 32); --Truncate to integer value
					
					extended_moved_y_bit_unsigned := moved_y * PIXEL_COEF; --Compute the pixel location
					truncated_extended_moved_y_bit_unsigned := extended_moved_y_bit_unsigned(32 + 9 downto 32); --Truncate to integer value
					inverted_y_bit := ROWS - truncated_extended_moved_y_bit_unsigned;
					moved_y_bit := std_logic_vector(inverted_y_bit);

					pixel_x <= moved_x_bit;
					pixel_y <= moved_y_bit;
					pixel_on <= "1";

					--Save the last rotated point and set current to be rotated
					if(point_position > 0) then
						rotated_points(point_position - 1).x := cordic_to_writer_x;
						rotated_points(point_position - 1).y := cordic_to_writer_y;
						unrotated_x <= points_to_draw(point_position).x;
						unrotated_y <= points_to_draw(point_position).y;
					end if;
					
					point_position := point_position + 1;

				else
					pixel_on <= "0";

					--Move the last point to the rotated points
					rotated_points(point_position - 1).x := cordic_to_writer_x;
					rotated_points(point_position - 1).y := cordic_to_writer_y;

					--Switch vectors
					points_to_draw := rotated_points;

				end if;



			end if;

		end if;

	end process;



end memory_writer_arq;