library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity Char_ROM is
	generic(
		N: integer:= 6;
		M: integer:= 3;
		W: integer:= 8
	);
	port(
		char_address: in std_logic_vector(5 downto 0);
		font_row, font_col: in std_logic_vector(M-1 downto 0);
		rom_out: out std_logic
	);
end;

architecture p of Char_ROM is
	subtype tipoLinea is std_logic_vector(0 to W-1);

	type char is array(0 to W-1) of tipoLinea;
	constant A: char:= (
								"00011000",
								"00111100",
								"01100110",
								"01100110",
								"01111110",
								"01100110",
								"01100110",
								"00000000"
						);
	constant B: char:= (
								"01111100",
								"01100110",
								"01100110",
								"01111100",
								"01100110",
								"01100110",
								"01111100",
								"00000000"
						);
	constant C: char:= (
								"00111110",
								"01100011",
								"01100000",
								"01100000",
								"01100000",
								"01100011",
								"00111110",
								"00000000"
						);

	constant D: char:= (
								"01111100",
								"01100110",
								"01100011",
								"01100011",
								"01100011",
								"01100110",
								"01111100",
								"00000000"
						);

	constant E: char:= (
								"01111110",
								"01100000",
								"01100000",
								"01111000",
								"01100000",
								"01100000",
								"01111110",
								"00000000"
						);

	constant F: char:= (
								"01111110",
								"01100000",
								"01100000",
								"01111000",
								"01100000",
								"01100000",
								"01100000",
								"00000000"
						);

	constant G: char:= (
								"00111100",
								"01100010",
								"01100000",
								"01101110",
								"01100110",
								"01100110",
								"00111100",
								"00000000"
						);

	constant H: char:= (
								"01100110",
								"01100110",
								"01100110",
								"01111110",
								"01100110",
								"01100110",
								"01100110",
								"00000000"
						);
						
	constant N_Char: char:= (
								"01100110",
								"01100110",
								"01110110",
								"01110110",
								"01101110",
								"01101110",
								"01100110",
								"00000000"
						);
						
	constant O: char:= ("00111100",
						"01111110",
						"11000111",
						"11001011",
						"11010011",
						"11100011",
						"01111110",
						"00111100"

						);


	constant ZERO: char:= (
						"00111100",
"01111110",
"11000111",
"11001011",
"11010011",
"11100011",
"01111110",
"00111100"
	
						);
	constant ONE: char:= (
						"00001000",
						"00011000",
						"00111000",
						"00011000",
						"00011000",
						"00011000",
						"01111110",
						"00000000");
						
	constant TWO: char:= (
	"00111100",
	"01100110",
	"01100110",
	"00001110",
	"00011100",
	"00111000",
	"01110110",
	"01111110"
);				
	constant THREE: char:= (
	"01111110",
	"01111110",
	"00000110",
	"01111110",
	"01111110",
	"00000110",
	"01111110",
	"01111110"
);				
	constant FOUR: char:= (
"00100110",
"01100110",
"01100110",
"01111110",
"00000110",
"00000110",
"00000110",
"00000110"
	
);				
	
	constant FIVE: char:= (
	
"01111110",
"01000110",
"01000000",
"01111100",
"01111110",
"00000010",
"01100010",
"01111110"
	
);				
	
	constant SIX: char:= (
	
"01111110",
"01000110",
"01000000",
"01000000",
"01111110",
"01100010",
"01100010",
"01111110"
	
	
);				
	
	
	constant SEVEN: char:= (
	
"01111110",
"01100010",
"00000110",
"00001100",
"00011000",
"00011000",
"00011000",
"00011000"
	
);				
	constant EIGHT: char:= (
"01111110",
"01000010",
"01000010",
"01000010",
"01111110",
"01000010",
"01000010",
"01111110"
	);				
	
	
	constant NINE: char:= (
"01111110",
"01100010",
"01100010",
"00111110",
"00011110",
"00000110",
"00000110",
"00000110"
);				
	
	constant COMMA: char:= (

"00000000",
"00000000",
"00000000",
"00000000",
"00011000",
"00011000",
"00001000",
"00010000"

	
	
	);
						
	constant Err: char:= (
								"00000000",
								"01111110",
								"01111110",
								"01100110",
								"01100110",
								"01111110",
								"01111110",
								"00000000"
						);
						
	constant SPACE: char:= (
								"00000000",
								"00000000",
								"00000000",
								"00000000",
								"00000000",
								"00000000",
								"00000000",
								"00000000"
						);
constant V: char:= (
								"11000011",
								"11000011",
								"01100110",
								"01100110",
								"00100100",
								"00011000",
								"00011000",
								"00000000"
						);										
	 

	type memo is array(0 to 255) of tipoLinea;
	signal RAM: memo:= (
								0 => ZERO(0), 1 => ZERO(1), 2 => ZERO(2), 3 => ZERO(3), 4 => ZERO(4), 5 => ZERO(5), 6 => ZERO(6), 7 => ZERO(7),
								8 => ONE(0), 9 => ONE(1), 10 => ONE(2), 11 => ONE(3), 12 => ONE(4), 13 => ONE(5), 14 => ONE(6), 15 => ONE(7),
								16 => TWO(0), 17 => TWO(1), 18 => TWO(2), 19 => TWO(3), 20 => TWO(4), 21 => TWO(5), 22 => TWO(6), 23 => TWO(7),
								24 => THREE(0), 25 => THREE(1), 26 => THREE(2), 27 => THREE(3), 28 => THREE(4), 29 => THREE(5), 30 => THREE(6), 31 => THREE(7),
								32 => FOUR(0), 33 => FOUR(1), 34 => FOUR(2), 35 => FOUR(3), 36 => FOUR(4), 37 => FOUR(5), 38 => FOUR(6), 39 => FOUR(7),
								40 => FIVE(0), 41 => FIVE(1), 42 => FIVE(2), 43 => FIVE(3), 44 => FIVE(4), 45 => FIVE(5), 46 => FIVE(6), 47 => FIVE(7),
								48 => SIX(0), 49 => SIX(1), 50 => SIX(2), 51 => SIX(3), 52 => SIX(4), 53 => SIX(5), 54 => SIX(6), 55 => SIX(7),
								56 => SEVEN(0), 57 => SEVEN(1), 58 => SEVEN(2), 59 => SEVEN(3), 60 => SEVEN(4), 61 => SEVEN(5), 62 => SEVEN(6), 63 => SEVEN(7),
								64 => EIGHT(0), 65 => EIGHT(1), 66 => EIGHT(2), 67 => EIGHT(3), 68 => EIGHT(4), 69 => EIGHT(5), 70 => EIGHT(6), 71 => EIGHT(7),
								72 => NINE(0), 73 => NINE(1), 74 => NINE(2), 75 => NINE(3), 76 => NINE(4), 77 => NINE(5), 78 => NINE(6), 79 => NINE(7),
								80 => COMMA(0), 81 => COMMA(1), 82 => COMMA(2), 83 => COMMA(3), 84 => COMMA(4), 85 => COMMA(5), 86 => COMMA(6), 87 => COMMA(7),
								88 => SPACE(0), 89 => SPACE(1), 90 => SPACE(2), 91 => SPACE(3), 92 => SPACE(4), 93 => SPACE(5), 94 => SPACE(6), 95 => SPACE(7),
								96 => V(0), 97 => V(1), 98 => V(2), 99 => V(3), 100 => V(4), 101 => V(5), 102 => V(6), 103 => V(7),
								104 to 255 => "00000000"
							);

	signal char_addr_aux: std_logic_vector(8 downto 0);
	
begin

	char_addr_aux <= char_address & font_row;
	rom_out <= RAM(conv_integer(char_addr_aux))(conv_integer(font_col));

end;