library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity Char_ROM is
	generic(
		N: integer:= 6;
		M: integer:= 3;
		W: integer:= 8
	);
	port(
		char_address: in std_logic_vector(5 downto 0);
		font_row, font_col: in std_logic_vector(M-1 downto 0);
		rom_out: out std_logic
	);
end;

architecture p of Char_ROM is
	subtype tipoLinea is std_logic_vector(0 to W-1);

	type char is array(0 to W-1) of tipoLinea;
	constant A: char:= (
								"00011000",
								"00111100",
								"01100110",
								"01100110",
								"01111110",
								"01100110",
								"01100110",
								"00000000"
						);
	constant B: char:= (
								"01111100",
								"01100110",
								"01100110",
								"01111100",
								"01100110",
								"01100110",
								"01111100",
								"00000000"
						);
	constant C: char:= (
								"00111110",
								"01100011",
								"01100000",
								"01100000",
								"01100000",
								"01100011",
								"00111110",
								"00000000"
						);

	constant D: char:= (
								"01111100",
								"01100110",
								"01100011",
								"01100011",
								"01100011",
								"01100110",
								"01111100",
								"00000000"
						);

	constant E: char:= (
								"01111110",
								"01100000",
								"01100000",
								"01111000",
								"01100000",
								"01100000",
								"01111110",
								"00000000"
						);

	constant F: char:= (
								"01111110",
								"01100000",
								"01100000",
								"01111000",
								"01100000",
								"01100000",
								"01100000",
								"00000000"
						);

	constant G: char:= (
								"00111100",
								"01100010",
								"01100000",
								"01101110",
								"01100110",
								"01100110",
								"00111100",
								"00000000"
						);

	constant H: char:= (
								"01100110",
								"01100110",
								"01100110",
								"01111110",
								"01100110",
								"01100110",
								"01100110",
								"00000000"
						);
						
	constant N_Char: char:= (
								"01100110",
								"01100110",
								"01110110",
								"01110110",
								"01101110",
								"01101110",
								"01100110",
								"00000000"
						);
						
	constant O: char:= (
								"00111100",
								"01100110",
								"01100110",
								"01100110",
								"01100110",
								"01100110",
								"00111100",
								"00000000"
						);
						
	constant Err: char:= (
								"00000000",
								"01111110",
								"01111110",
								"01100110",
								"01100110",
								"01111110",
								"01111110",
								"00000000"
						);
						

	type memo is array(0 to 255) of tipoLinea;
	signal RAM: memo:= (
								0 => A(0), 1 => A(1), 2 => A(2), 3 => A(3), 4 => A(4), 5 => A(5), 6 => A(6), 7 => A(7),
								8 => B(0), 9 => B(1), 10 => B(2), 11 => B(3), 12 => B(4), 13 => B(5), 14 => B(6), 15 => B(7),
								16 => C(0), 17 => C(1), 18 => C(2), 19 => C(3), 20 => C(4), 21 => C(5), 22 => C(6), 23 => C(7),
								24 => D(0), 25 => D(1), 26 => D(2), 27 => D(3), 28 => D(4), 29 => D(5), 30 => D(6), 31 => D(7),
								32 => E(0), 33 => E(1), 34 => E(2), 35 => E(3), 36 => E(4), 37 => E(5), 38 => E(6), 39 => E(7),
								40 => F(0), 41 => F(1), 42 => F(2), 43 => F(3), 44 => F(4), 45 => F(5), 46 => F(6), 47 => F(7),
								48 => G(0), 49 => G(1), 50 => G(2), 51 => G(3), 52 => G(4), 53 => G(5), 54 => G(6), 55 => G(7),
								56 => H(0), 57 => H(1), 58 => H(2), 59 => H(3), 60 => H(4), 61 => H(5), 62 => H(6), 63 => H(7),
								64 => N_Char(0), 65 => N_Char(1), 66 => N_Char(2), 67 => N_Char(3), 68 => N_Char(4), 69 => N_Char(5), 70 => N_Char(6), 71 => N_Char(7),
								72 => O(0), 73 => O(1), 74 => O(2), 75 => O(3), 76 => O(4), 77 => O(5), 78 => O(6), 79 => O(7),
								80 => Err(0), 81 => Err(1), 82 => Err(2), 83 => Err(3), 84 => Err(4), 85 => Err(5), 86 => Err(6), 87 => Err(7),
								88 to 255 => "00000000"
							);

	signal char_addr_aux: std_logic_vector(8 downto 0);
	
begin

	char_addr_aux <= char_address & font_row;
	rom_out <= RAM(conv_integer(char_addr_aux))(conv_integer(font_col));

end;