library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity tp1 is
  port (
		clk: in std_logic
	);
end;

architecture tp1_arq of tp1 is
begin

end;
